*KiCad schematic (cleaned for PSpice include)
.model D1 D
CBULK1 N_TVS1_K 0 10u
L1 N_TVS1_K INPUTSTAGEHV_BULK_P 1m
C1 INPUTSTAGEHV_BULK_P 0 10u
*TVS1 __TVS1
*J2 J2
Rf1 N_J1_Pin_1 N_F1_Pad1 10
D1 POWERVOUT_PLUS_INTERNAL POWERSW_NODE_INTERNAL __D1
CL1 POWERVOUT_PLUS_INTERNAL 0 330u
*U1 _U1
CVDD1 N_U1_VDD 0 100n
L2 POWERVOUT_PLUS_INTERNAL POWERSW_NODE_INTERNAL 1m
RFB1 FEEDBACKVOUT FEEDBACKFB_INTERNAL 10k
CFB1 FEEDBACKFB_INTERNAL 0 0.015u
RFB2 FEEDBACKFB_INTERNAL 0 121k