.title KiCad schematic
.model __D1 D
CBULK1 Net-_TVS1-K_ /POWER/VIN_MINUS 10U
L1 Net-_TVS1-K_ /INPUTSTAGE/HV_BULK_+ 2
C1 /INPUTSTAGE/HV_BULK_+ /POWER/VIN_MINUS 10U
TVS1 __TVS1
J2 __J2
Rf1 Net-_J1-Pin_1_ Net-_F1-Pad1_ 10
D1 /POWER/VOUT_PLUS_INTERNAL /POWER/SW_NODE_INTERNAL __D1
CL1 /POWER/VOUT_PLUS_INTERNAL /POWER/VIN_MINUS 330u
U1 __U1
CVDD1 Net-_U1-VDD_ /POWER/VIN_MINUS 100n
L2 /POWER/VOUT_PLUS_INTERNAL /POWER/SW_NODE_INTERNAL 1Meg
RFB1 /FEEDBACK/VOUT /FEEDBACK/FB_INTERNAL 10k
CFB1 /FEEDBACK/FB_INTERNAL /POWER/VIN_MINUS 0.015u
RFB2 /FEEDBACK/FB_INTERNAL /POWER/VIN_MINUS 121k
.end
