** Profile: "STARTUP-START_UP"  [ C:\Users\Oyebisi\Downloads\UCC28881 Stimulation files\UCC28881_PSPICE_TRANS\ucc28881_trans-pspicefiles\startup\start_up.sim ] 

** Creating circuit file "START_UP.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../ucc28881_trans.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 40n SKIPBP 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ITL1= 750
.OPTIONS ITL2= 100
.OPTIONS ITL4= 50
.OPTIONS RELTOL= 0.002
.PROBE64 V(alias(*)) I(alias(*)) 
.INC "..\STARTUP.net" 


.END
